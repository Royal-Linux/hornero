module hornero

pub const (
	version = '0.1.0'
)
